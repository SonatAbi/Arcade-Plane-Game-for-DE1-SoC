module waterpixel
    (input wire clk,
    input wire rst,
    input wire [10:0]  ox,
    input wire [10:0]  oy,
    input wire [10:0]  px,
    input wire [10:0]  py,
    output wire        water_color);

   wire 	             inobj;
   wire [6:0]  		 water_y, water_x;
	
   reg [31:0] 	       rom_data;
   wire [4:0] 	       rom_addr;
   wire               rom_bit;
	
   
   assign inobj     = (px >= ox) && (px < ox + 12'd128) && (py >=  oy) && (py < oy + 12'd128);
   
   assign water_x     = inobj ? px - ox : 0;
   assign water_y     = inobj ? py - oy : 0;
   
   assign rom_addr   = water_y[6:2];
   assign rom_bit    = rom_data[water_x[6:2]];
   
   assign water_color = (rom_bit) ? 1'b1 : 1'b0;

   always @*
     case (rom_addr)
       5'h00: rom_data = 32'b00000011000000000100000100000000; 
       5'h01: rom_data = 32'b00000100000000000100001000000011; 
       5'h02: rom_data = 32'b00001000000000001011101000011100; 
       5'h03: rom_data = 32'b00000100000000010000010001100000; 
       5'h04: rom_data = 32'b00001010000000100000010010010000; 
       5'h05: rom_data = 32'b00110010100001000000001010001110; 
       5'h06: rom_data = 32'b11000001010001000000001010000001; 
       5'h07: rom_data = 32'b00000010001010100000001001000000; 
       5'h08: rom_data = 32'b00000100000100010000110000100000; 
       5'h09: rom_data = 32'b00001000001000010001000000011000; 
       5'h0a: rom_data = 32'b11101000010000001010101010100100; 
       5'h0b: rom_data = 32'b00010100100000100100010001010011; 
       5'h0c: rom_data = 32'b00000101000001010000010001001100; 
       5'h0d: rom_data = 32'b00000011000001010000100001000001; 
       5'h0e: rom_data = 32'b00000001000001010000100010000001; 
       5'h0f: rom_data = 32'b11100000110010001001000100000010; 
       5'h10: rom_data = 32'b00011000001010001010001000000100; 
       5'h11: rom_data = 32'b00000100110001000100010111011000; 
       5'h12: rom_data = 32'b00000101000001000100010000100000; 
       5'h13: rom_data = 32'b00000010001101001100100001000000; 
       5'h14: rom_data = 32'b00000100010010010010100001000000; 
       5'h15: rom_data = 32'b00000100100010100001000001000000; 
       5'h16: rom_data = 32'b00011001000001000010000001000000; 
       5'h17: rom_data = 32'b11100010000001000100000010100000; 
       5'h18: rom_data = 32'b00010010000001010100000010001001; 
       5'h19: rom_data = 32'b00010001000010011000000100001010; 
       5'h1a: rom_data = 32'b11100000101100100100000010001010; 
       5'h1b: rom_data = 32'b00011000010000100010000100000100; 
       5'h1c: rom_data = 32'b00000101101000010001001000000100; 
       5'h1d: rom_data = 32'b00000010001000010000100100000100; 
       5'h1e: rom_data = 32'b00000001100100100000011011001000; 
       5'h1f: rom_data = 32'b00000000010101000000001000110000; 
     endcase
     
endmodule 